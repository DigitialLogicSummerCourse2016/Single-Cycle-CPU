`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr[30:2] < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin

ROMDATA[0] <= 32'b000010_00000_00000_00000_00000_000100; //RESET:  j INIT
ROMDATA[1] <= 32'b000010_00000_00000_00000_00001_101010; //ILLOP:  j INTRPT
ROMDATA[2] <= 32'b000010_00000_00000_00000_00000_000011; //XADR:  j EXPT
ROMDATA[3] <= 32'b000000_11111_00000_00000_00000_001000; //EXPT:  jr $ra
ROMDATA[4] <= 32'b000101_10001_00000_00000_00000_000100; //INIT:  bne $s1, $zero, START
ROMDATA[5] <= 32'b100011_11100_01000_00000_00000_001000; //   lw $t0, 8($gp)
ROMDATA[6] <= 32'b000101_01000_00000_00000_00000_000000; //   bne $t0, $zero, REPEAT
ROMDATA[7] <= 32'b001000_10001_10001_00000_00000_000001; //REPEAT:  addi $s1, $s1, 1
ROMDATA[8] <= 32'b000000_00000_00000_00000_00000_001000; //   jr $zero
ROMDATA[9] <= 32'b001000_00000_01000_00000_00000_111111; //START:  addi $t0, $zero, 0x3f
ROMDATA[10] <= 32'b101011_00000_01000_00000_00000_000000; // sw $t0, 0($zero)
ROMDATA[11] <= 32'b001000_00000_01001_00000_00000_000110; // addi $t1, $zero, 0x06
ROMDATA[12] <= 32'b101011_00000_01001_00000_00000_000100; // sw $t1, 4($zero)
ROMDATA[13] <= 32'b001000_00000_01000_00000_00001_011011; // addi $t0, $zero, 0x5b
ROMDATA[14] <= 32'b101011_00000_01000_00000_00000_001000; // sw $t0, 8($zero)
ROMDATA[15] <= 32'b001000_00000_01001_00000_00001_001111; // addi $t1, $zero, 0x4f
ROMDATA[16] <= 32'b101011_00000_01001_00000_00000_001100; // sw $t1, 12($zero)
ROMDATA[17] <= 32'b001000_00000_01000_00000_00001_100110; // addi $t0, $zero, 0x66
ROMDATA[18] <= 32'b101011_00000_01000_00000_00000_010000; // sw $t0, 16($zero)
ROMDATA[19] <= 32'b001000_00000_01001_00000_00001_101101; // addi $t1, $zero, 0x6d
ROMDATA[20] <= 32'b101011_00000_01001_00000_00000_010100; // sw $t1, 20($zero)
ROMDATA[21] <= 32'b001000_00000_01000_00000_00001_111101; // addi $t0, $zero, 0x7d
ROMDATA[22] <= 32'b101011_00000_01000_00000_00000_011000; // sw $t0, 24($zero)
ROMDATA[23] <= 32'b001000_00000_01001_00000_00000_000111; // addi $t1, $zero, 0x07
ROMDATA[24] <= 32'b101011_00000_01001_00000_00000_011100; // sw $t1, 28($zero)
ROMDATA[25] <= 32'b001000_00000_01000_00000_00001_111111; // addi $t0, $zero, 0x7f
ROMDATA[26] <= 32'b101011_00000_01000_00000_00000_100000; // sw $t0, 32($zero)
ROMDATA[27] <= 32'b001000_00000_01001_00000_00001_101111; // addi $t1, $zero, 0x6f
ROMDATA[28] <= 32'b101011_00000_01001_00000_00000_100100; // sw $t1, 36($zero)
ROMDATA[29] <= 32'b001000_00000_01000_00000_00001_110111; // addi $t0, $zero, 0x77
ROMDATA[30] <= 32'b101011_00000_01000_00000_00000_101000; // sw $t0, 40($zero)
ROMDATA[31] <= 32'b001000_00000_01001_00000_00001_111100; // addi $t1, $zero, 0x7c
ROMDATA[32] <= 32'b101011_00000_01001_00000_00000_101100; // sw $t1, 44($zero)
ROMDATA[33] <= 32'b001000_00000_01000_00000_00000_111001; // addi $t0, $zero, 0x39
ROMDATA[34] <= 32'b101011_00000_01000_00000_00000_110000; // sw $t0, 48($zero)
ROMDATA[35] <= 32'b001000_00000_01001_00000_00001_011110; // addi $t1, $zero, 0x5e
ROMDATA[36] <= 32'b101011_00000_01001_00000_00000_110100; // sw $t1, 52($zero)
ROMDATA[37] <= 32'b001000_00000_01000_00000_00001_111011; // addi $t0, $zero, 0x7b
ROMDATA[38] <= 32'b101011_00000_01000_00000_00000_111000; // sw $t0, 56($zero)
ROMDATA[39] <= 32'b001000_00000_01001_00000_00001_110001; // addi $t1, $zero, 0x71
ROMDATA[40] <= 32'b101011_00000_01001_00000_00000_111100; // sw $t1, 60($zero)
ROMDATA[41] <= 32'b001000_00000_10111_00000_00000_000001; // addi $s7, $zero, 1
ROMDATA[42] <= 32'b001111_00000_11100_01000_00000_000000; // lui $gp, 0x4000
ROMDATA[43] <= 32'b101011_11100_00000_00000_00000_001000; // sw $zero, 8($gp)
ROMDATA[44] <= 32'b001000_00000_01001_00000_00000_000011; // addi $t1, $zero, 3
ROMDATA[45] <= 32'b101011_11100_01001_00000_00000_100000; // sw $t1, 32($gp)
ROMDATA[46] <= 32'b001111_00000_01101_11111_11111_111111; // lui $t5, 0xffff
ROMDATA[47] <= 32'b001101_01101_01101_00111_10010_101111; // ori $t5, $t5, 0x3caf
ROMDATA[48] <= 32'b101011_11100_01101_00000_00000_000000; // sw $t5, 0($gp)
ROMDATA[49] <= 32'b101011_11100_01101_00000_00000_000100; // sw $t5, 4($gp)
ROMDATA[50] <= 32'b001000_00000_01110_00000_00000_000011; // addi $t6, $zero, 3
ROMDATA[51] <= 32'b101011_11100_01110_00000_00000_001000; // sw $t6, 8($gp)
ROMDATA[52] <= 32'b000010_00000_00000_00000_00000_110100; //STAY:  j STAY
ROMDATA[53] <= 32'b001000_11101_11101_11111_11111_110000; //bgcd:  addi $sp, $sp, -16
ROMDATA[54] <= 32'b101011_11101_10100_00000_00000_001100; // sw $s4, 12($sp)
ROMDATA[55] <= 32'b101011_11101_10010_00000_00000_001000; // sw $s2, 8($sp)
ROMDATA[56] <= 32'b101011_11101_10011_00000_00000_000100; // sw $s3, 4($sp)
ROMDATA[57] <= 32'b101011_11101_11111_00000_00000_000000; // sw $ra, 0($sp)
ROMDATA[58] <= 32'b000100_00100_00000_00000_00000_100001; // beq $a0, $zero, Return1
ROMDATA[59] <= 32'b000100_00101_00000_00000_00000_100010; // beq $a1, $zero, Return2
ROMDATA[60] <= 32'b001000_00000_01001_00000_00000_000001; // addi $t1, $zero, 1
ROMDATA[61] <= 32'b000000_00100_01001_10010_00000_100100; // and $s2, $a0, $t1
ROMDATA[62] <= 32'b000000_00101_01001_10011_00000_100100; // and $s3, $a1, $t1
ROMDATA[63] <= 32'b001000_00000_01001_00000_00000_000001; // addi $t1, $zero, 1
ROMDATA[64] <= 32'b000000_10010_10011_01010_00000_100101; // or $t2, $s2, $s3
ROMDATA[65] <= 32'b000101_01001_01010_00000_00000_000100; // bne $t1, $t2, ALLEVEN
ROMDATA[66] <= 32'b000000_10010_10011_01001_00000_100100; // and $t1, $s2, $s3
ROMDATA[67] <= 32'b000101_01001_00000_00000_00000_001100; // bne $t1, $zero, ALLODD
ROMDATA[68] <= 32'b000100_10010_00000_00000_00000_000101; // beq $s2, $zero, ONEEVEN
ROMDATA[69] <= 32'b000100_10011_00000_00000_00000_000111; // beq $s3, $zero, TWOEVEN
ROMDATA[70] <= 32'b000000_00000_00100_00100_00001_000010; //ALLEVEN: srl $a0, $a0, 1
ROMDATA[71] <= 32'b000000_00000_00101_00101_00001_000010; //     srl $a1, $a1, 1
ROMDATA[72] <= 32'b001000_10100_10100_00000_00000_000001; //     addi $s4, $s4, 1
ROMDATA[73] <= 32'b000011_00000_00000_00000_00000_110101; //     jal bgcd
ROMDATA[74] <= 32'b000000_00000_00100_00100_00001_000010; //ONEEVEN: srl $a0, $a0, 1
ROMDATA[75] <= 32'b000000_00101_00000_00101_00000_100000; // add $a1, $a1, $zero
ROMDATA[76] <= 32'b000011_00000_00000_00000_00000_110101; // jal bgcd
ROMDATA[77] <= 32'b000000_00000_00101_00101_00001_000010; //TWOEVEN: srl $a1, $a1, 1
ROMDATA[78] <= 32'b000000_00100_00000_00100_00000_100000; // add $a0, $a0, $zero
ROMDATA[79] <= 32'b000011_00000_00000_00000_00000_110101; // jal  bgcd
ROMDATA[80] <= 32'b000000_00100_00101_01001_00000_101010; //ALLODD:  slt $t1, $a0, $a1
ROMDATA[81] <= 32'b000101_01001_00000_00000_00000_000101; // bne $t1, $zero, ONELTWO
ROMDATA[82] <= 32'b000000_00100_00101_01001_00000_100010; // sub $t1, $a0, $a1
ROMDATA[83] <= 32'b000000_00000_01001_01001_00001_000010; // srl $t1, $t1, 1
ROMDATA[84] <= 32'b000000_01001_00000_00100_00000_100000; // add $a0 $t1, $zero
ROMDATA[85] <= 32'b000000_00101_00000_00101_00000_100000; // add $a1, $a1, $zero
ROMDATA[86] <= 32'b000011_00000_00000_00000_00000_110101; // jal bgcd
ROMDATA[87] <= 32'b000000_00101_00100_01001_00000_100010; //ONELTWO: sub $t1, $a1, $a0
ROMDATA[88] <= 32'b000000_00000_01001_01001_00001_000010; // srl $t1, $t1, 1
ROMDATA[89] <= 32'b000000_01001_00000_00101_00000_100000; // add $a1, $t1, $zero
ROMDATA[90] <= 32'b000000_00100_00000_00100_00000_100000; // add $a0, $a0, $zero
ROMDATA[91] <= 32'b000011_00000_00000_00000_00000_110101; // jal bgcd
ROMDATA[92] <= 32'b000000_00000_00101_00010_00000_100000; //Return1: add $v0, $zero, $a1
ROMDATA[93] <= 32'b000010_00000_00000_00000_00001_100000; // j LOOP
ROMDATA[94] <= 32'b000000_00000_00100_00010_00000_100000; //Return2: add $v0, $zero, $a0
ROMDATA[95] <= 32'b000010_00000_00000_00000_00001_100000; // j LOOP
ROMDATA[96] <= 32'b000100_10100_00000_00000_00000_000100; //LOOP:  beq $s4, $zero, GCDFIN
ROMDATA[97] <= 32'b000000_00000_00010_00010_00001_000000; // sll $v0, $v0, 1
ROMDATA[98] <= 32'b001000_00000_01001_00000_00000_000001; // addi $t1, $zero, 1
ROMDATA[99] <= 32'b000000_10100_01001_10100_00000_100010; // sub $s4, $s4, $t1
ROMDATA[100] <= 32'b000010_00000_00000_00000_00001_100000; // j LOOP
ROMDATA[101] <= 32'b101011_11100_00010_00000_00000_011000; //GCDFIN:  sw $v0, 24($gp)
ROMDATA[102] <= 32'b101011_11100_00010_00000_00000_001100; // sw $v0, 12($gp)
ROMDATA[103] <= 32'b001000_00000_01001_00000_00000_000011; // addi $t1, $zero, 3
ROMDATA[104] <= 32'b101011_11100_01001_00000_00000_100000; // sw $t1, 32($gp)
ROMDATA[105] <= 32'b000010_00000_00000_00000_00000_110100; // j STAY
ROMDATA[106] <= 32'b100011_11100_01111_00000_00000_100000; //INTRPT:  lw $t7, 32($gp)
ROMDATA[107] <= 32'b001010_01111_01001_00000_00000_001000; // slti $t1, $t7, 8
ROMDATA[108] <= 32'b000101_01001_00000_00000_00000_001110; // bne $t1, $zero, TIMER
ROMDATA[109] <= 32'b100011_11100_10000_00000_00000_011100; // lw $s0, 28($gp)
ROMDATA[110] <= 32'b000101_10110_00000_00000_00000_000100; // bne $s6, $zero, ALREADY
ROMDATA[111] <= 32'b000000_00000_10000_00100_00000_100000; // add $a0, $zero, $s0
ROMDATA[112] <= 32'b000000_00000_10000_11000_00000_100000; // add $t8, $zero, $s0
ROMDATA[113] <= 32'b001000_10110_10110_00000_00000_000001; // addi $s6, $s6, 1
ROMDATA[114] <= 32'b000000_11010_00000_00000_00000_001000; // jr $k0
ROMDATA[115] <= 32'b000000_00000_10000_00101_00000_100000; //ALREADY: add $a1, $zero, $s0
ROMDATA[116] <= 32'b000000_00000_10000_11001_00000_100000; // add $t9, $zero, $s0
ROMDATA[117] <= 32'b000000_00000_00000_10110_00000_100000; // add $s6, $zero, $zero
ROMDATA[118] <= 32'b000000_00000_00000_10000_00000_100000; // add $s0, $zero, $zero
ROMDATA[119] <= 32'b001000_00000_01001_00000_00000_000001; // addi $t1, $zero, 1
ROMDATA[120] <= 32'b101011_11100_01001_00000_00000_100000; // sw $t1, 32($gp)
ROMDATA[121] <= 32'b001000_11010_11010_00000_00000_000100; // addi $k0, $k0, 4
ROMDATA[122] <= 32'b000000_11010_00000_00000_00000_001000; // jr $k0
ROMDATA[123] <= 32'b001111_00000_01000_11111_11111_111111; //TIMER:  lui $t0, 0xffff
ROMDATA[124] <= 32'b001101_01000_01000_11111_11111_111001; // ori $t0, $t0, 0xfff9
ROMDATA[125] <= 32'b100011_11100_01001_00000_00000_001000; // lw $t1, 8($gp)
ROMDATA[126] <= 32'b000000_01001_01000_01001_00000_100100; // and $t1, $t1, $t0
ROMDATA[127] <= 32'b101011_11100_01001_00000_00000_001000; // sw $t1, 8($gp)
ROMDATA[128] <= 32'b000000_00000_10111_01010_01000_000000; //DIGI:  sll $t2, $s7, 8
ROMDATA[129] <= 32'b001010_01010_01111_00000_10000_000000; // slti $t7, $t2, 0x400
ROMDATA[130] <= 32'b000101_01111_00000_00000_00000_000111; // bne $t7, $zero, SECOND
ROMDATA[131] <= 32'b001010_01010_01110_00001_00000_000000; //FIRST:  slti $t6, $t2, 0x800
ROMDATA[132] <= 32'b000101_01110_00000_00000_00000_000011; // bne $t6, $zero FIRSTL
ROMDATA[133] <= 32'b001100_11000_01100_00000_00011_110000; //FIRSTH:  andi $t4, $t8, 0x00f0
ROMDATA[134] <= 32'b000000_00000_01100_01100_00100_000010; // srl $t4, $t4, 4
ROMDATA[135] <= 32'b000010_00000_00000_00000_00010_010000; // j DISPLAY
ROMDATA[136] <= 32'b001100_11000_01100_00000_00000_001111; //FIRSTL:  andi $t4, $t8, 0x000f
ROMDATA[137] <= 32'b000010_00000_00000_00000_00010_010000; // j DISPLAY
ROMDATA[138] <= 32'b001010_01010_01110_00000_01000_000000; //SECOND:  slti  $t6, $t2, 0x200
ROMDATA[139] <= 32'b000101_01110_00000_00000_00000_000011; // bne $t6, $zero, SECONDL
ROMDATA[140] <= 32'b001100_11001_01100_00000_00011_110000; //SECONDH: andi $t4, $t9, 0x00f0
ROMDATA[141] <= 32'b000000_00000_01100_01100_00100_000010; // srl $t4, $t4, 4
ROMDATA[142] <= 32'b000010_00000_00000_00000_00010_010000; // j DISPLAY
ROMDATA[143] <= 32'b001100_11001_01100_00000_00000_001111; //SECONDL: andi $t4, $t9, 0x000f
ROMDATA[144] <= 32'b000000_00000_01100_01100_00010_000000; //DISPLAY: sll $t4, $t4, 2
ROMDATA[145] <= 32'b100011_01100_01100_00000_00000_000000; // lw $t4, 0($t4)
ROMDATA[146] <= 32'b000000_01010_01100_01010_00000_100000; // add $t2, $t2, $t4
ROMDATA[147] <= 32'b101011_11100_01010_00000_00000_010100; // sw $t2, 20($gp)
ROMDATA[148] <= 32'b000000_00000_10111_10111_00001_000000; // sll $s7, $s7, 1
ROMDATA[149] <= 32'b001010_10111_01110_00000_00000_001001; // slti $t6, $s7, 0x09
ROMDATA[150] <= 32'b000101_01110_00000_00000_00000_000001; // bne $t6, $zero, FIN
ROMDATA[151] <= 32'b001000_00000_10111_00000_00000_000001; // addi $s7, $zero, 1
ROMDATA[152] <= 32'b100011_11100_01001_00000_00000_001000; //FIN:  lw $t1, 8($gp)
ROMDATA[153] <= 32'b001101_01001_01001_00000_00000_000010; // ori $t1, $t1, 0x0002
ROMDATA[154] <= 32'b101011_11100_01001_00000_00000_001000; // sw $t1, 8($gp)
ROMDATA[155] <= 32'b000000_11010_00000_00000_00000_001000; // jr $k0
//no error

		for (i=156;i<ROM_SIZE;i=i+1) begin
			ROMDATA[i] <= 32'b0;
		end
end
endmodule
