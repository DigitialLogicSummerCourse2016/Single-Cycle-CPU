`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 128;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr[30:2] < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin

//		ROMDATA[0] <= 32'h3c094000;
//		ROMDATA[1] <= 32'h3525001c;
//		ROMDATA[2] <= 32'h8ca20000;
//		ROMDATA[3] <= 32'h00023020;
//		ROMDATA[4] <= 32'h8ca20000;
//		ROMDATA[5] <= 32'h00023820;
//		ROMDATA[6] <= 32'h00c78820;
//		ROMDATA[7] <= 32'hacb1fffc;

//		ROMDATA[0] <= 32'h3c114000;
//		ROMDATA[1] <= 32'h26310004;
//		ROMDATA[2] <= 32'h241000aa;
//		ROMDATA[3] <= 32'hae200000;
//		ROMDATA[4] <= 32'h08100000;
//		ROMDATA[5] <= 32'h0c000000;
//		ROMDATA[6] <= 32'h00000000;
//		ROMDATA[7] <= 32'h3402000a;
//		ROMDATA[8] <= 32'h0000000c;
//		ROMDATA[9] <= 32'h0000_0000;
//		ROMDATA[10]<= 32'h0274_8825;
//		ROMDATA[11] <= 32'h0800_0015;
//		ROMDATA[12] <= 32'h0274_8820;
//		ROMDATA[13] <= 32'h0800_0015;
//		ROMDATA[14] <= 32'h0274_882A;
//		ROMDATA[15] <= 32'h1011_0002;
//		ROMDATA[16] <= 32'h0293_8822;
//		ROMDATA[17] <= 32'h0800_0015;
//		ROMDATA[18] <= 32'h0274_8822;
//		ROMDATA[19] <= 32'h0800_0015;
//		ROMDATA[20] <= 32'h0274_8824;
//		ROMDATA[21] <= 32'hae11_0003;
//		ROMDATA[22] <= 32'h0800_0001;
//
//	    for (i=23;i<ROM_SIZE;i=i+1) begin
//            ROMDATA[i] <= 32'b0;
//        end

			ROMDATA[0] <= 32'b00001000000100000000000000000100;
			ROMDATA[1] <= 32'b00001000000100000000000001100010;
			ROMDATA[2] <= 32'b00001000000100000000000000000011;
			ROMDATA[3] <= 32'b00000011111000000000000000001000;
			ROMDATA[4] <= 32'b00100000000010000000000000111111;
			ROMDATA[5] <= 32'b10101100000010000000000000000000;
			ROMDATA[6] <= 32'b00100000000010010000000000000110;
			ROMDATA[7] <= 32'b10101100000010010000000000000100;
			ROMDATA[8] <= 32'b00100000000010000000000001011011;
			ROMDATA[9] <= 32'b10101100000010000000000000001000;
			ROMDATA[10] <= 32'b00100000000010010000000001001111;
			ROMDATA[11] <= 32'b10101100000010010000000000001100;
			ROMDATA[12] <= 32'b00100000000010000000000001100110;
			ROMDATA[13] <= 32'b10101100000010000000000000010000;
			ROMDATA[14] <= 32'b00100000000010010000000001101101;
			ROMDATA[15] <= 32'b10101100000010010000000000010100;
			ROMDATA[16] <= 32'b00100000000010000000000001111101;
			ROMDATA[17] <= 32'b10101100000010000000000000011000;
			ROMDATA[18] <= 32'b00100000000010010000000000000111;
			ROMDATA[19] <= 32'b10101100000010010000000000011100;
			ROMDATA[20] <= 32'b00100000000010000000000001111111;
			ROMDATA[21] <= 32'b10101100000010000000000000100000;
			ROMDATA[22] <= 32'b00100000000010010000000001101111;
			ROMDATA[23] <= 32'b10101100000010010000000000100100;
			ROMDATA[24] <= 32'b00100000000010000000000001110111;
			ROMDATA[25] <= 32'b10101100000010000000000000101000;
			ROMDATA[26] <= 32'b00100000000010010000000001111100;
			ROMDATA[27] <= 32'b10101100000010010000000000101100;
			ROMDATA[28] <= 32'b00100000000010000000000000111001;
			ROMDATA[29] <= 32'b10101100000010000000000000110000;
			ROMDATA[30] <= 32'b00100000000010010000000001011110;
			ROMDATA[31] <= 32'b10101100000010010000000000110100;
			ROMDATA[32] <= 32'b00100000000010000000000001111011;
			ROMDATA[33] <= 32'b10101100000010000000000000111000;
			ROMDATA[34] <= 32'b00100000000010010000000001110001;
			ROMDATA[35] <= 32'b10101100000010010000000000111100;
			ROMDATA[36] <= 32'b00100000000101110000000000000001;
			ROMDATA[37] <= 32'b00000000000000001011100000100000;
			ROMDATA[38] <= 32'b00111100000111000100000000000000;
			ROMDATA[39] <= 32'b10101111101000000000000000001000;
			ROMDATA[40] <= 32'b00100000000010010000000000000011;
			ROMDATA[41] <= 32'b10101111100010010000000000100000;
			ROMDATA[42] <= 32'b00001000000100000000000000101010;
			ROMDATA[43] <= 32'b00111100000011011111111111111110;
			ROMDATA[44] <= 32'b00110101101011010111100101011111;
			ROMDATA[45] <= 32'b10101111100011010000000000000000;
			ROMDATA[46] <= 32'b00110101101011011111111111111111;
			ROMDATA[47] <= 32'b10101111100011010000000000000100;
			ROMDATA[48] <= 32'b00100000000011100000000000000011;
			ROMDATA[49] <= 32'b10101111100011100000000000001000;
			ROMDATA[50] <= 32'b00100011101111011111111111110000;
			ROMDATA[51] <= 32'b10101111101101000000000000001100;
			ROMDATA[52] <= 32'b10101111101100100000000000001000;
			ROMDATA[53] <= 32'b10101111101100110000000000000100;
			ROMDATA[54] <= 32'b10101111101111110000000000000000;
			ROMDATA[55] <= 32'b00010000100000000000000000100001;
			ROMDATA[56] <= 32'b00010000101000000000000000100010;
			ROMDATA[57] <= 32'b00100000000010010000000000000001;
			ROMDATA[58] <= 32'b00000000100010011001000000100100;
			ROMDATA[59] <= 32'b00000000101010011001100000100100;
			ROMDATA[60] <= 32'b00100000000010010000000000000001;
			ROMDATA[61] <= 32'b00000010010100110101000000100101;
			ROMDATA[62] <= 32'b00010101001010100000000000000100;
			ROMDATA[63] <= 32'b00000010010100110100100000100100;
			ROMDATA[64] <= 32'b00010101001000000000000000001100;
			ROMDATA[65] <= 32'b00010010010000000000000000000101;
			ROMDATA[66] <= 32'b00010010011000000000000000000111;
			ROMDATA[67] <= 32'b00000000000001000010000001000010;
			ROMDATA[68] <= 32'b00000000000001010010100001000010;
			ROMDATA[69] <= 32'b00100010100101000000000000000001;
			ROMDATA[70] <= 32'b00001100000100000000000000110010;
			ROMDATA[71] <= 32'b00000000000001000010000001000010;
			ROMDATA[72] <= 32'b00000000101000000010100000100000;
			ROMDATA[73] <= 32'b00001100000100000000000000110010;
			ROMDATA[74] <= 32'b00000000000001010010100001000010;
			ROMDATA[75] <= 32'b00000000100000000010000000100000;
			ROMDATA[76] <= 32'b00001100000100000000000000110010;
			ROMDATA[77] <= 32'b00000000100001010100100000101010;
			ROMDATA[78] <= 32'b00010101001000000000000000000101;
			ROMDATA[79] <= 32'b00000000100001010100100000100010;
			ROMDATA[80] <= 32'b00000000000010010100100001000010;
			ROMDATA[81] <= 32'b00000001001000000010000000100000;
			ROMDATA[82] <= 32'b00000000101000000010100000100000;
			ROMDATA[83] <= 32'b00001100000100000000000000110010;
			ROMDATA[84] <= 32'b00000000101001000100100000100010;
			ROMDATA[85] <= 32'b00000000000010010100100001000010;
			ROMDATA[86] <= 32'b00000001001000000010100000100000;
			ROMDATA[87] <= 32'b00000000100000000010000000100000;
			ROMDATA[88] <= 32'b00001100000100000000000000110010;
			ROMDATA[89] <= 32'b00000000000001010001000000100000;
			ROMDATA[90] <= 32'b00001000000100000000000001011101;
			ROMDATA[91] <= 32'b00000000000001000001000000100000;
			ROMDATA[92] <= 32'b00001000000100000000000001011101;
			ROMDATA[93] <= 32'b00010010100000001111111111001100;
			ROMDATA[94] <= 32'b00000000000000100001000001000000;
			ROMDATA[95] <= 32'b00100000000010010000000000000001;
			ROMDATA[96] <= 32'b00000010100010011010000000100010;
			ROMDATA[97] <= 32'b00001000000100000000000001011101;
			ROMDATA[98] <= 32'b10001111100011110000000000100000;
			ROMDATA[99] <= 32'b00101001111010010000000000001000;
			ROMDATA[100] <= 32'b00010101001000000000000000001010;
			ROMDATA[101] <= 32'b10001111100000110000000000011100;
			ROMDATA[102] <= 32'b00010110110000000000000000000011;
			ROMDATA[103] <= 32'b00000000000000110010000000100000;
			ROMDATA[104] <= 32'b00100010110101100000000000000001;
			ROMDATA[105] <= 32'b00000011010000000000000000001000;
			ROMDATA[106] <= 32'b00000000000000110010100000100000;
			ROMDATA[107] <= 32'b00000000000000001011000000100000;
			ROMDATA[108] <= 32'b00000000000000000001100000100000;
			ROMDATA[109] <= 32'b00100011010110100000000000000100;
			ROMDATA[110] <= 32'b00000011010000000000000000001000;
			ROMDATA[111] <= 32'b00111100000010001111111111111111;
			ROMDATA[112] <= 32'b00110101000010001111111111111001;
			ROMDATA[113] <= 32'b10001111100010010000000000001000;
			ROMDATA[114] <= 32'b00000001001010000100100000100100;
			ROMDATA[115] <= 32'b10101111100010010000000000001000;
			ROMDATA[116] <= 32'b00010100010000000000000000000001;
			ROMDATA[117] <= 32'b10101111100000100000000000001100;
			ROMDATA[118] <= 32'b00000000000101110101001000000000;
			ROMDATA[119] <= 32'b00101001010011110000010000000000;
			ROMDATA[120] <= 32'b00010101111000000000000000000111;
			ROMDATA[121] <= 32'b00101001010011100000100000000000;
			ROMDATA[122] <= 32'b00010101110000000000000000000011;
			ROMDATA[123] <= 32'b00110000100011000000000011110000;
			ROMDATA[124] <= 32'b00000000000011000110000100000010;
			ROMDATA[125] <= 32'b00001000000100000000000010000110;
			ROMDATA[126] <= 32'b00110000100011000000000000001111;
			ROMDATA[127] <= 32'b00001000000100000000000010000110;
			ROMDATA[128] <= 32'b00101001010011100000001000000000;
			ROMDATA[129] <= 32'b00010101110000000000000000000011;
			ROMDATA[130] <= 32'b00110000101011000000000011110000;
			ROMDATA[131] <= 32'b00000000000011000110000100000010;
			ROMDATA[132] <= 32'b00001000000100000000000010000110;
			ROMDATA[133] <= 32'b00110000101011000000000000001111;
			ROMDATA[134] <= 32'b00000000000011000110000010000000;
			ROMDATA[135] <= 32'b10001101100011000000000000000000;
			ROMDATA[136] <= 32'b00000001010011000101000000100000;
			ROMDATA[137] <= 32'b10101111101010100000000000010100;
			ROMDATA[138] <= 32'b00000000000101111011100001000000;
			ROMDATA[139] <= 32'b00101010111011100000000000001001;
			ROMDATA[140] <= 32'b00010101110000000000000000000001;
			ROMDATA[141] <= 32'b00100000000101110000000000000001;
			ROMDATA[142] <= 32'b10001111100010010000000000001000;
			ROMDATA[143] <= 32'b00110101001010010000000000000010;
			ROMDATA[144] <= 32'b10101111100010010000000000001000;
			ROMDATA[145] <= 32'b00000011010000000000000000001000;


		for (i=146;i<ROM_SIZE;i=i+1) begin
			ROMDATA[i] <= 32'b0;
		end
end
endmodule
