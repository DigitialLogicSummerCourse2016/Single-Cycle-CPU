`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 128;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr[30:2] < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin

//			ROMDATA[0] <= 32'b00001000000100000000000000000100;
//			ROMDATA[1] <= 32'b00001000000100000000000001100010;
//			ROMDATA[2] <= 32'b00001000000100000000000000000011;
//			ROMDATA[3] <= 32'b00000011111000000000000000001000;
//			ROMDATA[4] <= 32'b00100000000010000000000000111111;
//			ROMDATA[5] <= 32'b10101100000010000000000000000000;
//			ROMDATA[6] <= 32'b00100000000010010000000000000110;
//			ROMDATA[7] <= 32'b10101100000010010000000000000100;
//			ROMDATA[8] <= 32'b00100000000010000000000001011011;
//			ROMDATA[9] <= 32'b10101100000010000000000000001000;
//			ROMDATA[10] <= 32'b00100000000010010000000001001111;
//			ROMDATA[11] <= 32'b10101100000010010000000000001100;
//			ROMDATA[12] <= 32'b00100000000010000000000001100110;
//			ROMDATA[13] <= 32'b10101100000010000000000000010000;
//			ROMDATA[14] <= 32'b00100000000010010000000001101101;
//			ROMDATA[15] <= 32'b10101100000010010000000000010100;
//			ROMDATA[16] <= 32'b00100000000010000000000001111101;
//			ROMDATA[17] <= 32'b10101100000010000000000000011000;
//			ROMDATA[18] <= 32'b00100000000010010000000000000111;
//			ROMDATA[19] <= 32'b10101100000010010000000000011100;
//			ROMDATA[20] <= 32'b00100000000010000000000001111111;
//			ROMDATA[21] <= 32'b10101100000010000000000000100000;
//			ROMDATA[22] <= 32'b00100000000010010000000001101111;
//			ROMDATA[23] <= 32'b10101100000010010000000000100100;
//			ROMDATA[24] <= 32'b00100000000010000000000001110111;
//			ROMDATA[25] <= 32'b10101100000010000000000000101000;
//			ROMDATA[26] <= 32'b00100000000010010000000001111100;
//			ROMDATA[27] <= 32'b10101100000010010000000000101100;
//			ROMDATA[28] <= 32'b00100000000010000000000000111001;
//			ROMDATA[29] <= 32'b10101100000010000000000000110000;
//			ROMDATA[30] <= 32'b00100000000010010000000001011110;
//			ROMDATA[31] <= 32'b10101100000010010000000000110100;
//			ROMDATA[32] <= 32'b00100000000010000000000001111011;
//			ROMDATA[33] <= 32'b10101100000010000000000000111000;
//			ROMDATA[34] <= 32'b00100000000010010000000001110001;
//			ROMDATA[35] <= 32'b10101100000010010000000000111100;
//			ROMDATA[36] <= 32'b00100000000101110000000000000001;
//			ROMDATA[37] <= 32'b00000000000000001011100000100000;
//			ROMDATA[38] <= 32'b00111100000111000100000000000000;
//			ROMDATA[39] <= 32'b10101111101000000000000000001000;
//			ROMDATA[40] <= 32'b00100000000010010000000000000011;
//			ROMDATA[41] <= 32'b10101111100010010000000000100000;
//			ROMDATA[42] <= 32'b00001000000100000000000000101010;
//			ROMDATA[43] <= 32'b00111100000011011111111111111110;
//			ROMDATA[44] <= 32'b00110101101011010111100101011111;
//			ROMDATA[45] <= 32'b10101111100011010000000000000000;
//			ROMDATA[46] <= 32'b00110101101011011111111111111111;
//			ROMDATA[47] <= 32'b10101111100011010000000000000100;
//			ROMDATA[48] <= 32'b00100000000011100000000000000011;
//			ROMDATA[49] <= 32'b10101111100011100000000000001000;
//			ROMDATA[50] <= 32'b00100011101111011111111111110000;
//			ROMDATA[51] <= 32'b10101111101101000000000000001100;
//			ROMDATA[52] <= 32'b10101111101100100000000000001000;
//			ROMDATA[53] <= 32'b10101111101100110000000000000100;
//			ROMDATA[54] <= 32'b10101111101111110000000000000000;
//			ROMDATA[55] <= 32'b00010000100000000000000000100001;
//			ROMDATA[56] <= 32'b00010000101000000000000000100010;
//			ROMDATA[57] <= 32'b00100000000010010000000000000001;
//			ROMDATA[58] <= 32'b00000000100010011001000000100100;
//			ROMDATA[59] <= 32'b00000000101010011001100000100100;
//			ROMDATA[60] <= 32'b00100000000010010000000000000001;
//			ROMDATA[61] <= 32'b00000010010100110101000000100101;
//			ROMDATA[62] <= 32'b00010101001010100000000000000100;
//			ROMDATA[63] <= 32'b00000010010100110100100000100100;
//			ROMDATA[64] <= 32'b00010101001000000000000000001100;
//			ROMDATA[65] <= 32'b00010010010000000000000000000101;
//			ROMDATA[66] <= 32'b00010010011000000000000000000111;
//			ROMDATA[67] <= 32'b00000000000001000010000001000010;
//			ROMDATA[68] <= 32'b00000000000001010010100001000010;
//			ROMDATA[69] <= 32'b00100010100101000000000000000001;
//			ROMDATA[70] <= 32'b00001100000100000000000000110010;
//			ROMDATA[71] <= 32'b00000000000001000010000001000010;
//			ROMDATA[72] <= 32'b00000000101000000010100000100000;
//			ROMDATA[73] <= 32'b00001100000100000000000000110010;
//			ROMDATA[74] <= 32'b00000000000001010010100001000010;
//			ROMDATA[75] <= 32'b00000000100000000010000000100000;
//			ROMDATA[76] <= 32'b00001100000100000000000000110010;
//			ROMDATA[77] <= 32'b00000000100001010100100000101010;
//			ROMDATA[78] <= 32'b00010101001000000000000000000101;
//			ROMDATA[79] <= 32'b00000000100001010100100000100010;
//			ROMDATA[80] <= 32'b00000000000010010100100001000010;
//			ROMDATA[81] <= 32'b00000001001000000010000000100000;
//			ROMDATA[82] <= 32'b00000000101000000010100000100000;
//			ROMDATA[83] <= 32'b00001100000100000000000000110010;
//			ROMDATA[84] <= 32'b00000000101001000100100000100010;
//			ROMDATA[85] <= 32'b00000000000010010100100001000010;
//			ROMDATA[86] <= 32'b00000001001000000010100000100000;
//			ROMDATA[87] <= 32'b00000000100000000010000000100000;
//			ROMDATA[88] <= 32'b00001100000100000000000000110010;
//			ROMDATA[89] <= 32'b00000000000001010001000000100000;
//			ROMDATA[90] <= 32'b00001000000100000000000001011101;
//			ROMDATA[91] <= 32'b00000000000001000001000000100000;
//			ROMDATA[92] <= 32'b00001000000100000000000001011101;
//			ROMDATA[93] <= 32'b00010010100000001111111111001100;
//			ROMDATA[94] <= 32'b00000000000000100001000001000000;
//			ROMDATA[95] <= 32'b00100000000010010000000000000001;
//			ROMDATA[96] <= 32'b00000010100010011010000000100010;
//			ROMDATA[97] <= 32'b00001000000100000000000001011101;
//			ROMDATA[98] <= 32'b10001111100011110000000000100000;
//			ROMDATA[99] <= 32'b00101001111010010000000000001000;
//			ROMDATA[100] <= 32'b00010101001000000000000000001010;
//			ROMDATA[101] <= 32'b10001111100000110000000000011100;
//			ROMDATA[102] <= 32'b00010110110000000000000000000011;
//			ROMDATA[103] <= 32'b00000000000000110010000000100000;
//			ROMDATA[104] <= 32'b00100010110101100000000000000001;
//			ROMDATA[105] <= 32'b00000011010000000000000000001000;
//			ROMDATA[106] <= 32'b00000000000000110010100000100000;
//			ROMDATA[107] <= 32'b00000000000000001011000000100000;
//			ROMDATA[108] <= 32'b00000000000000000001100000100000;
//			ROMDATA[109] <= 32'b00100011010110100000000000000100;
//			ROMDATA[110] <= 32'b00000011010000000000000000001000;
//			ROMDATA[111] <= 32'b00111100000010001111111111111111;
//			ROMDATA[112] <= 32'b00110101000010001111111111111001;
//			ROMDATA[113] <= 32'b10001111100010010000000000001000;
//			ROMDATA[114] <= 32'b00000001001010000100100000100100;
//			ROMDATA[115] <= 32'b10101111100010010000000000001000;
//			ROMDATA[116] <= 32'b00010100010000000000000000000001;
//			ROMDATA[117] <= 32'b10101111100000100000000000001100;
//			ROMDATA[118] <= 32'b00000000000101110101001000000000;
//			ROMDATA[119] <= 32'b00101001010011110000010000000000;
//			ROMDATA[120] <= 32'b00010101111000000000000000000111;
//			ROMDATA[121] <= 32'b00101001010011100000100000000000;
//			ROMDATA[122] <= 32'b00010101110000000000000000000011;
//			ROMDATA[123] <= 32'b00110000100011000000000011110000;
//			ROMDATA[124] <= 32'b00000000000011000110000100000010;
//			ROMDATA[125] <= 32'b00001000000100000000000010000110;
//			ROMDATA[126] <= 32'b00110000100011000000000000001111;
//			ROMDATA[127] <= 32'b00001000000100000000000010000110;
//			ROMDATA[128] <= 32'b00101001010011100000001000000000;
//			ROMDATA[129] <= 32'b00010101110000000000000000000011;
//			ROMDATA[130] <= 32'b00110000101011000000000011110000;
//			ROMDATA[131] <= 32'b00000000000011000110000100000010;
//			ROMDATA[132] <= 32'b00001000000100000000000010000110;
//			ROMDATA[133] <= 32'b00110000101011000000000000001111;
//			ROMDATA[134] <= 32'b00000000000011000110000010000000;
//			ROMDATA[135] <= 32'b10001101100011000000000000000000;
//			ROMDATA[136] <= 32'b00000001010011000101000000100000;
//			ROMDATA[137] <= 32'b10101111101010100000000000010100;
//			ROMDATA[138] <= 32'b00000000000101111011100001000000;
//			ROMDATA[139] <= 32'b00101010111011100000000000001001;
//			ROMDATA[140] <= 32'b00010101110000000000000000000001;
//			ROMDATA[141] <= 32'b00100000000101110000000000000001;
//			ROMDATA[142] <= 32'b10001111100010010000000000001000;
//			ROMDATA[143] <= 32'b00110101001010010000000000000010;
//			ROMDATA[144] <= 32'b10101111100010010000000000001000;
//			ROMDATA[145] <= 32'b00000011010000000000000000001000;

			ROMDATA[0] <= 32'b00001000000000000000000000000011; //Start: j    Reset
			ROMDATA[1] <= 32'b00001000000000000000000001000110; //ILLOP: j    Intrpt
			ROMDATA[2] <= 32'b00001000000000000000000001000101; //XADR: j    Expt
			ROMDATA[3] <= 32'b00000000000000001110100000100000; //Reset: add  $sp  , $0  , $0
			ROMDATA[4] <= 32'b00100000000010000000000011111100; // addi $t0  , $0  , 0xfc
			ROMDATA[5] <= 32'b10101111101010000000000000000000; // sw   $t0  , 0($sp)
			ROMDATA[6] <= 32'b00100000000010010000000001100000; // addi $t1  , $0  , 0x60
			ROMDATA[7] <= 32'b10101111101010010000000000000100; // sw   $t1  , 4 ($sp)
			ROMDATA[8] <= 32'b00100000000010000000000011011010; // addi $t0  , $0  , 0xda
			ROMDATA[9] <= 32'b10101111101010000000000000001000; // sw   $t0  , 8 ($sp)
			ROMDATA[10] <= 32'b00100000000010010000000011110010; // addi $t1  , $0  , 0xf2
			ROMDATA[11] <= 32'b10101111101010010000000000001100; // sw   $t1  , 12($sp)
			ROMDATA[12] <= 32'b00100000000010000000000001100110; // addi $t0  , $0  , 0x66
			ROMDATA[13] <= 32'b10101111101010000000000000010000; // sw   $t0  , 16($sp)
			ROMDATA[14] <= 32'b00100000000010010000000010110110; // addi $t1  , $0  , 0xb6
			ROMDATA[15] <= 32'b10101111101010010000000000010100; // sw   $t1  , 20($sp)
			ROMDATA[16] <= 32'b00100000000010000000000010111110; // addi $t0  , $0  , 0xbe
			ROMDATA[17] <= 32'b10101111101010000000000000011000; // sw   $t0  , 24($sp)
			ROMDATA[18] <= 32'b00100000000010010000000011100000; // addi $t1  , $0  , 0xe0
			ROMDATA[19] <= 32'b10101111101010010000000000011100; // sw   $t1  , 28($sp)
			ROMDATA[20] <= 32'b00100000000010000000000011111110; // addi $t0  , $0  , 0xfe
			ROMDATA[21] <= 32'b10101111101010000000000000100000; // sw   $t0  , 32($sp)
			ROMDATA[22] <= 32'b00100000000010010000000011110110; //    addi $t1  , $0  , 0xf6
			ROMDATA[23] <= 32'b10101111101010010000000000100100; // sw   $t1  , 36($sp)
			ROMDATA[24] <= 32'b00100000000010000000000011101110; // addi $t0  , $0  , 0xee
			ROMDATA[25] <= 32'b10101111101010000000000000101000; // sw   $t0  , 40($sp)
			ROMDATA[26] <= 32'b00100000000010010000000000111110; // addi $t1  , $0  , 0x3e
			ROMDATA[27] <= 32'b10101111101010010000000000101100; // sw   $t1  , 44($sp)
			ROMDATA[28] <= 32'b00100000000010000000000010011100; // addi $t0  , $0  , 0x9c
			ROMDATA[29] <= 32'b10101111101010000000000000110000; // sw   $t0  , 48($sp)
			ROMDATA[30] <= 32'b00100000000010010000000001111010; // addi $t1  , $0  , 0x7a
			ROMDATA[31] <= 32'b10101111101010010000000000110100; // sw   $t1  , 52($sp)
			ROMDATA[32] <= 32'b00100000000010000000000010011110; // addi $t0  , $0  , 0x9e
			ROMDATA[33] <= 32'b10101111101010000000000000111000; // sw   $t0  , 56($sp)
			ROMDATA[34] <= 32'b00100000000010010000000010001110; // addi $t1  , $0  , 0x8e
			ROMDATA[35] <= 32'b10101111101010010000000000111100; // sw   $t1  , 60($sp)
			ROMDATA[36] <= 32'b00100000000101100000000000000001; // addi $s6  , $0  , 1
			ROMDATA[37] <= 32'b00000000000000001011100000100000; // add  $s7  , $0  , $0
			ROMDATA[38] <= 32'b00111100000011010100000000000000; // lui  $t5  , 0x00004000
			ROMDATA[39] <= 32'b00110101101111010000000000000000; // ori  $sp  , $t5 , 0x00000000
			ROMDATA[40] <= 32'b00100000000010010000000000000011; // addi $t1  , $0  , 3
			ROMDATA[41] <= 32'b10101111101010010000000000100000; // sw   $t1  , 32($sp)
			ROMDATA[42] <= 32'b10101111101000000000000000001000; // sw   $0   , 8 ($sp)
			ROMDATA[43] <= 32'b00000000000000001110100000100000; // add  $sp  , $0  , $0
			ROMDATA[44] <= 32'b00001000000000000000000000101100; //Read: j    Read
			ROMDATA[45] <= 32'b00111100000011010100000000000000; //main: lui  $t5  , 0x00004000
			ROMDATA[46] <= 32'b00110101101111010000000000000000; // ori  $sp  , $t5 , 0x00000000
			ROMDATA[47] <= 32'b00111100000011011111111111111111; // lui  $t5  , 0xffff
			ROMDATA[48] <= 32'b00110100000100011111111100000000; // ori  $s1  , $0  , 0xff00
			ROMDATA[49] <= 32'b00000010001011011000100000100000; // add  $s1  , $s1 , $t5
			ROMDATA[50] <= 32'b10101111101100010000000000000000; // sw   $s1  , 0($sp)
			ROMDATA[51] <= 32'b10101111101100010000000000000100; // sw   $s1  , 4($sp)
			ROMDATA[52] <= 32'b00100000000100100000000000000011; // addi $s2  , $0  , 3
			ROMDATA[53] <= 32'b10101111101100100000000000001000; // sw   $s2  , 8($sp)
			ROMDATA[54] <= 32'b00000010100000000010000000100000; // add  $a0  , $s4 , $0
			ROMDATA[55] <= 32'b00000010101000000010100000100000; // add  $a1  , $s5 , $0
			ROMDATA[56] <= 32'b00000000000000000001000000100000; // add  $v0  , $0  , $0
			ROMDATA[57] <= 32'b00010000100001010000000000000111; //GCD: beq  $a0  , $a1 , Result
			ROMDATA[58] <= 32'b00000000100001010001100000100010; // sub  $v1  , $a0 , $a1
			ROMDATA[59] <= 32'b00000000011000000001100000101010; // slt  $v1  , $v1 , $0
			ROMDATA[60] <= 32'b00010000011000000000000000000010; // beq  $v1  , $0  , A
			ROMDATA[61] <= 32'b00000000101001000010100000100010; // sub  $a1  , $a1 , $a0
			ROMDATA[62] <= 32'b00001000000000000000000000111001; // j    GCD
			ROMDATA[63] <= 32'b00000000100001010010000000100010; //A: sub  $a0  , $a0 , $a1
			ROMDATA[64] <= 32'b00001000000000000000000000111001; // j    GCD
			ROMDATA[65] <= 32'b00000000100001010010000000100010; //Result: sub  $a0  , $a0 , $a1
			ROMDATA[66] <= 32'b10101111101001010000000000011000; // sw   $a1  , 24($sp)
			ROMDATA[67] <= 32'b00000000000000001110100000100000; // add  $sp  , $0  , $0
			ROMDATA[68] <= 32'b00001000000000000000000000101100; // j    Read
			ROMDATA[69] <= 32'b00000011111000000000000000001000; //Expt: jr   $ra
			ROMDATA[70] <= 32'b00000011101000000100000000100000; //Intrpt: add  $t0  , $sp ,$0
			ROMDATA[71] <= 32'b00111100000000010100000000000000; // lui  $at  , 0x00004000
			ROMDATA[72] <= 32'b00110100001111010000000000000000; // ori  $sp  , $at , 0x00000000
			ROMDATA[73] <= 32'b10001111101100110000000000100000; // lw   $s3  , 32($sp)
			ROMDATA[74] <= 32'b00101010011011110000000000001000; // slti $t7  , $s3 , 8
			ROMDATA[75] <= 32'b00010101111000000000000000001101; // bne  $t7  , $0  , Timer
			ROMDATA[76] <= 32'b10001111101000100000000000011100; //UART: lw   $v0  , 28($sp)
			ROMDATA[77] <= 32'b00010110111000000000000000000100; // bne  $s7  , $0  , Save2
			ROMDATA[78] <= 32'b00000000010000001010000000100000; //Save1: add  $s4  , $v0 , $0
			ROMDATA[79] <= 32'b00100010111101110000000000000001; // addi $s7  , $s7 , 1
			ROMDATA[80] <= 32'b00000001000000001110100000100000; // add  $sp  , $t0 , $0
			ROMDATA[81] <= 32'b00000011010000000000000000001000; // jr   $k0
			ROMDATA[82] <= 32'b00000000000000001011100000100000; //Save2: add  $s7  , $0  , $0
			ROMDATA[83] <= 32'b00000000010000001010100000100000; // add  $s5  , $v0 , $0
			ROMDATA[84] <= 32'b00100000000010010000000000000001; // addi $t1  , $0  , 1
			ROMDATA[85] <= 32'b10101111101010010000000000100000; // sw   $t1  , 32($sp)
			ROMDATA[86] <= 32'b00000001000000001110100000100000; // add  $sp  , $t0 , $0
			ROMDATA[87] <= 32'b00100011010110100000000000000100; // addi $k0  , $k0 , 4
			ROMDATA[88] <= 32'b00000011010000000000000000001000; // jr   $k0
			ROMDATA[89] <= 32'b00111100000000011111111111111111; //Timer: lui  $at  , 0x0000ffff
			ROMDATA[90] <= 32'b00110100001000011111111111111001; // ori  $at  , $at , 0x0000fff9
			ROMDATA[91] <= 32'b00000010010000011001000000100100; // and  $s2  , $s2 , $at
			ROMDATA[92] <= 32'b10101111101100100000000000001000; // sw   $s2  , 8 ($sp)
			ROMDATA[93] <= 32'b00010100100000000000000000000001; // bne  $a0  , $0  , DIGI
			ROMDATA[94] <= 32'b10101111101001010000000000001100; //LEDS: sw   $a1  , 12($sp)
			ROMDATA[95] <= 32'b00000000000101100111001000000000; //DIGI: sll  $t6  , $s6 , 8
			ROMDATA[96] <= 32'b00101001110011110000010000000000; // slti $t7  , $t6 , 0x400
			ROMDATA[97] <= 32'b00010101111000000000000000000111; // bne  $t7  , $0  , Load2
			ROMDATA[98] <= 32'b00101001110011110000100000000000; //Load1:     slti $t7  , $t6 , 0x800
			ROMDATA[99] <= 32'b00010001111000000000000000000010; // beq  $t7  , $0  , Load1H
			ROMDATA[100] <= 32'b00110010100011000000000000001111; //Load1L: andi $t4  , $s4 , 0x000f
			ROMDATA[101] <= 32'b00001000000000000000000001101000; // j    Load1Fin
			ROMDATA[102] <= 32'b00110010100011000000000011110000; //Load1H: andi $t4  , $s4 , 0x00f0
			ROMDATA[103] <= 32'b00000000000011000110000100000010; // srl  $t4  , $t4 , 4
			ROMDATA[104] <= 32'b00001000000000000000000001101111; //Load1Fin:     j    Display
			ROMDATA[105] <= 32'b00101001110011110000001000000000; //Load2: slti $t7  , $t6 , 0x200
			ROMDATA[106] <= 32'b00010001111000000000000000000010; // beq  $t7  , $0  , Load2H
			ROMDATA[107] <= 32'b00110010101011000000000000001111; //Load2L: andi $t4  , $s5 , 0x000f
			ROMDATA[108] <= 32'b00001000000000000000000001101111; // j    Display
			ROMDATA[109] <= 32'b00110010101011000000000011110000; //Load2H: andi $t4  , $s5 , 0x00f0
			ROMDATA[110] <= 32'b00000000000011000110000100000010; // srl  $t4  , $t4 , 4
			ROMDATA[111] <= 32'b00000000000011000110000010000000; //Display: sll  $t4  , $t4 , 2
			ROMDATA[112] <= 32'b10001101100011000000000000000000; //    lw   $t4  , 0 ($t4)
			ROMDATA[113] <= 32'b00000001110011000111000000100000; // add  $t6  , $t6 , $t4
			ROMDATA[114] <= 32'b10101111101011100000000000010100; // sw   $t6  , 20($sp)
			ROMDATA[115] <= 32'b00000000000101101011000001000000; // sll  $s6  , $s6 , 1
			ROMDATA[116] <= 32'b00101010110011100000000000001001; // slti $t6  , $s6 , 9
			ROMDATA[117] <= 32'b00010101110000000000000000000001; // bne  $t6  , $0  , Intrpt_Fin
			ROMDATA[118] <= 32'b00100000000101100000000000000001; // addi $s6  , $0  , 1
			ROMDATA[119] <= 32'b00110110010100100000000000000010; //Intrpt_Fin: ori  $s2  , $s2 , 0x00000002
			ROMDATA[120] <= 32'b10101111101100100000000000001000; // sw   $s2  , 8 ($sp)
			ROMDATA[121] <= 32'b00000001000000001110100000100000; // add  $sp  , $t0 , $0
			ROMDATA[122] <= 32'b00000011010000000000000000001000; // jr   $k0

		for (i=123;i<ROM_SIZE;i=i+1) begin
			ROMDATA[i] <= 32'b0;
		end

//		for (i=146;i<ROM_SIZE;i=i+1) begin
//			ROMDATA[i] <= 32'b0;
//		end
end
endmodule
